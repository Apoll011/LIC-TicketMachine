LIBRARY ieee;
USE ieee.std_logic_1164.all;

entity TicketMachine is
	port(
		RESET, CLK  	: in std_logic
	);
end TicketMachine;

architecture logicFunction OF TicketMachine IS
begin

END logicFunction;